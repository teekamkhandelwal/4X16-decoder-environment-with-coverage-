///PACKET
`ifndef _base_
`define _base_
class pkt;
  randc bit [3:0] x;
 rand bit e;
bit [15:0] d;
endclass
`endif
