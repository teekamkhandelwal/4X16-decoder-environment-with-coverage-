//TOP
`include "pkt.sv"
`include "interface.sv"
`include "gen.sv"
`include "driver.sv"
`include "monitor.sv"
`include "sb.sv"
`include "env.sv"
module top();
df_intf intf();
decoder d2(intf);
env e1(intf);
endmodule
